-- Testbench for mclk_gen module
