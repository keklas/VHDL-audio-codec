library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity mclk_gen is
    port (
        
    );
end mclk_gen;

architecture rtl of mclk_gen is

begin

end architecture;
