-- Testbench for ac_audio module