library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity ac_audio is
    port (
        
    );
end ac_audio;

architecture rtl of ac_audio is

begin

end architecture;