library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity ac_control is
    port (
        
    );
end ac_control;

architecture rtl of ac_control is

begin

end architecture;