-- Testbench for ac_control module